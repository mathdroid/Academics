-- PRAKTIKUM EL 3111 ARSITEKTUR SISTEM KOMPUTER
-- MODUL 4
-- PERCOBAAN 2
-- 17 NOV 2014
-- KELOMPOK VI
-- ROMBONGAN A
-- DAMON PRASETYO ARSO (13212001)
-- MUHAMMAD MUSTADI (13210056)
-- leftshift.vhdl
-- PROGRAM PENGGESER 2 BIT
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
LIBRARY altera_mf;
USE altera_mf.altera_mf_components.ALL;


ENTITY lshift_32_32 IS
  PORT (
    D_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0); -- Input 32-bit;
    D_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0) -- Output 32-bit;
    );
END lshift_32_32;ENTITY lshift_26_28 ISPORT (D_IN : IN STD_LOGIC_VECTOR (25 DOWNTO 0); -- Input 26-bit;D_OUT : OUT STD_LOGIC_VECTOR (27 DOWNTO 0) -- Output 28-bit;);END lshift_26_28;ARCHITECTURE behavior OF lshift_32_32 IS  BEGIN  D_OUT(31 DOWNTO 2) <= D_IN(29 DOWNTO 0);  D_OUT(1 DOWNTO 0) <= "00";END behavior;ARCHITECTURE behavior OF lshift_26_28 IS  BEGIN  D_OUT(27 DOWNTO 2) <= D_IN(25 DOWNTO 0);  D_OUT(1 DOWNTO 0) <= "00";END behavior;