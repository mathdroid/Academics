-- PRAKTIKUM EL 3111 ARSITEKTUR SISTEM KOMPUTER
-- MODUL 4
-- PERCOBAAN 2
-- 17 NOV 2014
-- KELOMPOK VI
-- ROMBONGAN A
-- DAMON PRASETYO ARSO (13212001)
-- MUHAMMAD MUSTADI (13210056)
-- cla32.vhdl
-- CARRY LOOK ADDER
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
LIBRARY altera_mf;
USE altera_mf.altera_mf_components.ALL;

ENTITY ALU IS
PORT (
  OPRND_1 : IN std_logic_vector (31 DOWNTO 0); -- Data Input 1
  OPRND_2 : IN std_logic_vector (31 DOWNTO 0); -- Data Input 2
  OP_SEL : IN std_logic; -- Operation Select
  RESULT : OUT std_logic_vector (31 DOWNTO 0) -- Data Output
);
END ALU;

ARCHITECTURE structure OF ALU IS
  COMPONENT cla32
    PORT (
      OPRND_1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      OPRND_2 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      C_IN : IN STD_LOGIC;
      RESULT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      C_OUT : OUT STD_LOGIC
      );
  END COMPONENT;
  FOR ALL : cla32 USE ENTITY cla_32(behavior);
  BEGIN
    cla32_1 : cla32 PORT MAP(OPRND_1=>OPRND_1, OPRND_2=>OPRND_2,C_IN=>OP_SEL,RESULT=>RESULT);
END structure;
